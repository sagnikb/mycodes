Shunt Clipper DC analysis
r1 1 2 1k
*default diode p-n
d1 2 3
*independent DC source - 2V
vdc 3 0 dc 2
*independent DC source with varying voltage
vin 1 0 dc 0
*DC analysis on source vin, to vary from -5V to +5V
.dc vin -5 5 0.01
.control
run
plot v(2) vs v(1)
.endc
.end
